`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:33:04 10/03/2016 
// Design Name: 
// Module Name:    top_module 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module top_module(
	output idle_LED
   );	
	 
	wire [10:0] href, vref;
	wire buffer_read, image_sel;
	
	dual_image_buffer imgbuf(
		.href, // from microblaze, 0-751
		.vref, // 0-480
		.fifo_data, // 8 bit data in from fifo
		.fifo_rck, // 1MHz clock signal generated by FPGA
		.get_data(buffer_read), // enable a new read sequence
		.image_sel(image_sel),
		.buffer_ready, // indicate that buffer has been filled
		.fifo_rrst, // fifo read reset (reset read addr pointer to 0)
		.fifo_oe, // fifo output enable (allow for addr pointer to increment)
		.pixel_value, // 8-bit value from internal buffer
		.trigger
   );

	disparity disp(
		.clk, // Read clk signal
		.enable, // enable new disparity calculation 
		.reset, // reset disparity FSM
		.image_data, // FIFO data in
		.buffer_ready,
		.new_image(buffer_read),
		.buffer_href,
		.buffer_vref,
		.image_sel(image_sel), // left/right frame select
		.idle(idle_LED) // LED indicator signify end of process
    );
	
	endmodule
