`timescale 1ns / 1ps

module ZedCamTest_top(
    input sysclk,
    input reset, // reset 
    input cam_rst, // button for camera RESET_BAR
    input trigger, // button for camera trigger
    input SW_camSelect, // switch for camera output enable
    input SW_read_fifo,
    output cam_sysclk, // sysclk out to camera
    output cam_reset, // reset_bar out to camera
    output cam_trigger, // trigger out to camera
    output i2c_ready, // LED indicator for i2c bus ready
    input output_sel,
    input [10:0] xLoc,
    input [10:0] yLoc,
    output [7:0] pixel_out,
    input [7:0] FIFO_DATA, // DO[7:0] from AL422b fifo
    output FIFO_OE1, // read enable to fifo (active low)
    output FIFO_RRST1, // read reset to fifo (active low)
    output FIFO_OE2, // read enable to fifo (active low)
    output FIFO_RRST2, // read reset to fifo (active low)
    output FIFO_RCK, // rck to fifo (1MHz)
    output [7:0] rgb, // values on vga color pins
    output HS, // horizontal sync (to VGA port)
    output VS // vertical sync (to VGA port)
);
    
wire clk_20Hz, clk_10kHz, clk_1MHz, clk_5MHz, clk_24MHz, clk_25MHz;

clk_wiz_0 mmcm(// Clock in ports
      .clk_in1(sysclk),
      // Clock out ports
      .clk_out1(clk_25MHz),
      .clk_out2(clk_24MHz),
      .clk_out3(clk_5MHz)
     );
     
// further divide the dcm clock to other freqs	 
clk_divs clks(
      .reset(reset), // synchronous reset
      .clk_24M(clk_24MHz), // 24MHz camera SCLK
      .clk_fifo(clk_1MHz), // 1MHz FIFO RCK
      .clk_debounce(clk_20Hz), // 20Hz clock pulse for debouncing stuff
      .anodes(clk_10kHz) // 10k 7Seg anode driver
     );
     
assign cam_sysclk = clk_24MHz;
assign FIFO_RCK = clk_5MHz;

// camera initialization sequence
reg [11:0] init_count = 12'h000;
always @(posedge clk_24MHz) // cam sysclk before ODDR2
begin
	if (cam_rst) // if cam_rst is pressed, redo the initialization sequence
	begin
		init_count <= 12'h000;
	end
	else if(init_count < 2500) // keep cam_rst asserted for at least 20 cam_sysclk cycles - I use 30 since it's the minimum time for the i2c bus to be ready
		init_count <= init_count + 1'b1;
end
assign cam_reset = (init_count >= 20);
assign i2c_ready = (init_count >= 30);

wire read_en;
debounce fifoRead_en(
    .clk(clk_20Hz),
    .btn(SW_read_fifo),
    .btn_val(read_en)
    );

wire cam_sel;
debounce camSelector(
    .clk(clk_20Hz),
    .btn(SW_camSelect),
    .btn_val(cam_sel)
    );

wire get_data;
debounce trig(
    .clk(clk_20Hz),
    .btn(trigger),
    .btn_val(get_data)
    );

wire fifo_rden, fifo_read_en, fifo_reset; //also connected to fifo_buffer
assign FIFO_OE1 = cam_sel == 1'b0 ? fifo_rden : 1'b1;
assign FIFO_RRST1 = cam_sel == 1'b0 ? fifo_reset : 1'b1;
assign FIFO_OE2 = cam_sel == 1'b1 ? fifo_rden : 1'b1;
assign FIFO_RRST2 = cam_sel == 1'b1 ? fifo_reset : 1'b1;

wire [7:0] pixelVal; // value of a camera pixel from fpga line buffer -> microblaze
wire [10:0] hc,hcount; // pixel number on current line
wire [10:0] vc,vcount; // number of current line
wire blank;

vga_controller_640_60 vgaOut(
	.rst(reset), 
	.pixel_clk(clk_25MHz),
	.HS(HS),
	.VS(VS),
	.hcount(hcount),
	.vcount(vcount),
	.blank(blank) 
);

assign hc = output_sel == 1'b0 ? hcount : xLoc;
assign vc = output_sel == 1'b0 ? vcount : yLoc;
assign rgb = output_sel == 1'b0 ? pixelVal : 8'h00;
assign pixel_out = output_sel == 1'b0 ? 8'h00 : pixelVal;

imgbuf fifo_buffer(
    .get_data(get_data),
	.href(hc),
	.vref(vc),
	.blank(blank),
	.fifo_data(FIFO_DATA), // 8 bit data in from fifo
	.fifo_rck(clk_5MHz), // 1MHz clock signal generated by FPGA
	.vga_clk(clk_25MHz),
	.fifo_rrst(fifo_reset), // fifo read reset (reset read addr pointer to 0)
	.fifo_oe(fifo_rden), // fifo output enable (allow for addr pointer to increment)
	.pixel_value(pixelVal), // 8-bit pixel value from internal buffer
	//.current_line(),
	.trigger(cam_trigger)
   );
   
endmodule
