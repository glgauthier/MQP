`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module for reading from the AL422b FIFO and storing pixel line data in a 
// local buffer.
//////////////////////////////////////////////////////////////////////////////////
module dual_image_buffer(
	input [10:0] href, // from microblaze, 0-751
	input [10:0] vref, // 0-480
	input [7:0] fifo_data, // 8 bit data in from fifo
	input fifo_rck, // 1MHz clock signal generated by FPGA
	input reg get_data, // enable a new read sequence
	input image_sel, // left/right image data out
   output reg buffer_ready, // indicate that buffer has been filled
	output reg fifo_rrst, // fifo read reset (reset read addr pointer to 0)
	output reg fifo_oe, // fifo output enable (allow for addr pointer to increment)
	output reg [7:0] pixel_value, // 8-bit value from internal buffer
	output reg trigger
   );

reg reset_pointer; 

parameter [1:0] ready = 2'b00;
parameter [1:0] read = 2'b01;
parameter [1:0] done = 2'b10;  
parameter [1:0] init = 2'b11;
reg buffer_ready;

reg [1:0] state = ready;
reg [1:0] prev_state, next_state = ready;

reg [7:0] pixel_array [0:59][0:91]; // implemented in BRAM

reg [9:0] pixel = 10'b00_0000_0000;
reg [15:0] num_lines = 16'h0000;

always @(posedge fifo_rck)
	state <= next_state;
	
always @(state,get_data,num_lines,pixel)	
	case(state)
		ready: 
			begin
				if(get_data) 
				begin
					trigger = 1'b0;
					next_state = init;
				end
				else
					next_state = ready;
					
				prev_state = ready;
			end
		init: 
			begin
				next_state = read;
				prev_state = init;
			end
		read: 
			begin
				if(num_lines == 280) // was pixel == 751
					next_state = done;
				else
					next_state = read;
					
				prev_state = read;
			end
		done: 
			begin
				next_state = ready;
				prev_state = done;
				trigger = 1'b1;
			end
	endcase

always @(posedge fifo_rck)
begin
		if(state==ready) // allow for MCS to read from pixel_line
			begin
			fifo_rrst <= 1'b1; // make sure read addr doesn't get reset
			end
		else if(state == init) // prepare to read new data from the AL422 into pixel_line
			begin
			pixel <= 10'b00_0000_000;
			buffer_ready <= 1'b0;
			fifo_oe <= 1'b0; // allow for read pointer to increment
			end
		else if(state == read) // read data in from the AL422
			begin
			if(next_state == done)
				fifo_oe <= 1'b1; // turn off read enable
			
			if((prev_state != init) && (pixel < 751)) // one cycle delay between init and valid data
				
				if((pixel>=329 && pixel <= 421) && (num_lines >= 209 && num_lines <= 269)) // read in top left corner of image
				begin
					pixel_array[(num_lines-209)][(pixel-329)] <= fifo_data;
					pixel <= pixel + 1'b1;
				end
				else
					pixel <= pixel + 1'b1;
			else if(prev_state != init)
				begin
				pixel <= 10'b00_0000_0000;
				num_lines <= num_lines + 1'b1;
				end
			end
		else if(state == done)
			begin
			buffer_ready <= 1'b1;
			fifo_rrst <= 1'b0;
			num_lines <= 16'h0000;
			end
end

// allow for input to read stored pixel line at given addr if state==ready
always @ (href, vref, pixel_value, pixel_array)
	pixel_value [7:0] = pixel_array[vref][href];



endmodule